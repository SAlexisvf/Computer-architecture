library IEEE;use IEEE.STD_LOGIC_1164.ALL;use IEEE.NUMERIC_STD.ALL;library UNISIM;use UNISIM.VComponents.all;
entity ROM is	PORT(		DIRECCION : IN STD_LOGIC_VECTOR(31 DOWNTO 0);		DATO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)	);end ROM;
architecture Behavioral of ROM isbegin
PROCESS(DIRECCION)
SUBTYPE REGISTRO IS STD_LOGIC_VECTOR(31 DOWNTO 0);TYPE REG_BANK IS ARRAY(0 TO 31) OF REGISTRO; 
VARIABLE ROM_MEMORY : REG_BANK := ( 
	x"0001_0004",	x"0002_0003",	x"0003_0002",	x"0004_0001",
	x"1111_1111",OTHERS => (OTHERS => '0') );BEGIN	DATO <= ROM_MEMORY(TO_INTEGER(UNSIGNED(DIRECCION(6 downto 2))));END PROCESS;
end Behavioral;

